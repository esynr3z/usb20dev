//==============================================================================
// Package with global types and parameters
//
//------------------------------------------------------------------------------
// 2018, Eden Synrez <esynr3z@gmail.com>
//==============================================================================

package usb_pkg;

typedef logic [7:0]  bus8_t;
typedef logic [31:0] bus32_t;

endpackage : usb_pkg
