//==============================================================================
// Package with global types and parameters
//
//------------------------------------------------------------------------------
// [usb20dev] 2018 Eden Synrez <esynr3z@gmail.com>
//==============================================================================

package usb_pkg;

parameter STUFF_BITS_N = 6;

typedef logic [7:0]  bus8_t;
typedef logic [31:0] bus32_t;

endpackage : usb_pkg
